`define LW_CMD 			0
`define PS_CMD 			1
`define PSI_CMD 		2
//-------------------------------------------------------
`define ADD_CMD 		8
`define ADDI_CMD 		9
`define MUL_CMD 		10
`define MULI_CMD 		11
`define SUB_CMD 		12
`define SUBI_CMD 		13
`define DIV_CMD 		14
`define DIVI_CMD 		15
//--------------------------------------------------------
`define OR_CMD 			16
`define ORI_CMD 		17
`define AND_CMD 		18
`define ANDI_CMD 		19
`define XOR_CMD 		20
`define XORI_CMD 		21
`define INV_CMD 		22
//--------------------------------------------------------
`define J_CMD 			24
`define JAL_CMD 		25
`define JR_CMD 			26
`define JL_CMD 			27
//--------------------------------------------------------
`define SLL_CMD 		32
`define SLLV_CMD 		33
`define SRL_CMD 		34
`define SRLV_CMD 		35
`define SLA_CMD 		36
`define SRA_CMD 		37
//--------------------------------------------------------
`define BEQ_CMD 		40
`define BQE_CMD 		41
`define BGERAL_CMD 	42
`define BGTZ_CMD 		43
`define BLEZ_CMD 		44
`define BLTZ_CMD 		45
`define BNE_CMD 		46